module RAM16K(out,en,clk,address,in,rw);
input[15:0]in;
input[13:0]address;
input rw,en,clk;
output[15:0]out;
wire en0,en1,en2,en3,msb13,msb12;
wire[11:0]rest0;
wire[15:0]out0,out1,out2,out3,out4,out5;
BUFFER buff0(msb13,address[13]);
BUFFER buff1(msb12,address[12]);
BUFFER buff2(rest0[11],address[11]);
BUFFER buff3(rest0[10],address[10]);
BUFFER buff4(rest0[9],address[9]);
BUFFER buff5(rest0[8],address[8]);
BUFFER buff6(rest0[7],address[7]);
BUFFER buff7(rest0[6],address[6]);
BUFFER buff8(rest0[5],address[5]);
BUFFER buff9(rest0[4],address[4]);
BUFFER buff10(rest0[3],address[3]);
BUFFER buff11(rest0[2],address[2]);
BUFFER buff12(rest0[1],address[1]);
BUFFER buff13(rest0[0],address[0]);
DEMUX_4WAY demux1(en0,en1,en2,en3,msb13,msb12,en);
RAM4K ram1(out0,en0,clk,rest0,in,rw);
RAM4K ram2(out1,en1,clk,rest0,in,rw);
RAM4K ram3(out2,en2,clk,rest0,in,rw);
RAM4K ram4(out3,en3,clk,rest0,in,rw);
OR_16_BIT_GATE or1(out4,out0,out1);
OR_16_BIT_GATE or2(out5,out2,out4);
OR_16_BIT_GATE or3(out,out3,out5);
endmodule
