module RAM4K(out,en,clk,address,in,rw);
input[15:0]in;
input[11:0]address;
input rw,en,clk;
output[15:0]out;
wire msb11,msb10,msb9,en0,en1,en2,en3,en4,en5,en6,en7;
wire[8:0]rest0;
wire[15:0]out0,out1,out2,out3,out4,out5,out6,out7,out8,out9,out10,out11,out12,out13;
BUFFER buff1(msb11,address[11]);
BUFFER buff2(msb10,address[10]);
BUFFER buff3(msb9,address[9]);
BUFFER buff4(rest0[8],address[8]);
BUFFER buff5(rest0[7],address[7]);
BUFFER buff6(rest0[6],address[6]);
BUFFER buff7(rest0[5],address[5]);
BUFFER buff8(rest0[4],address[4]);
BUFFER buff9(rest0[3],address[3]);
BUFFER buff10(rest0[2],address[2]);
BUFFER buff11(rest0[1],address[1]);
BUFFER buff12(rest0[0],address[0]);
DEMUX_8WAY demux1(en0,en1,en2,en3,en4,en5,en6,en7,msb9,msb10,msb11,en);
RAM512 ram1(out0,en0,clk,rest0,in,rw);
RAM512 ram2(out1,en1,clk,rest0,in,rw);
RAM512 ram3(out2,en2,clk,rest0,in,rw);
RAM512 ram4(out3,en3,clk,rest0,in,rw);
RAM512 ram5(out4,en4,clk,rest0,in,rw);
RAM512 ram6(out5,en5,clk,rest0,in,rw);
RAM512 ram7(out6,en6,clk,rest0,in,rw);
RAM512 ram8(out7,en7,clk,rest0,in,rw);
OR_16_BIT_GATE or1(out8,out0,out1);
OR_16_BIT_GATE or2(out9,out2,out8);
OR_16_BIT_GATE or3(out10,out3,out9);
OR_16_BIT_GATE or4(out11,out4,out10);
OR_16_BIT_GATE or5(out12,out5,out11);
OR_16_BIT_GATE or6(out13,out6,out12);
OR_16_BIT_GATE or7(out,out7,out13);
endmodule
